module Inverse_Mix_Columns(
    input CLK,
    input [0:127] INPUT,
    output [0:127] OUTPUT
    );

wire [0:31] Column_1, Column_2, Column_3, Column_4;

wire [0:7] C11, C12, C13, C14;
wire [0:7] C21, C22, C23, C24;
wire [0:7] C31, C32, C33, C34;
wire [0:7] C41, C42, C43, C44;

wire [0:7] Q10, Q11, Q12, Q13, Q14, Q15, Q16, Q17, Q18, Q19, Q110, Q111, Q112, Q113, Q114, Q115;
wire [0:7] Q20, Q21, Q22, Q23, Q24, Q25, Q26, Q27, Q28, Q29, Q210, Q211, Q212, Q213, Q214, Q215;
wire [0:7] Q30, Q31, Q32, Q33, Q34, Q35, Q36, Q37, Q38, Q39, Q310, Q311, Q312, Q313, Q314, Q315;
wire [0:7] Q40, Q41, Q42, Q43, Q44, Q45, Q46, Q47, Q48, Q49, Q410, Q411, Q412, Q413, Q414, Q415;

assign Column_1 = INPUT[0:31];
assign Column_2 = INPUT[32:63];
assign Column_3 = INPUT[64:95];
assign Column_4 = INPUT[96:127];

assign C11 = Column_1[0:7];
assign C12 = Column_1[8:15];
assign C13 = Column_1[16:23];
assign C14 = Column_1[24:31];

assign C21 = Column_2[0:7];
assign C22 = Column_2[8:15];
assign C23 = Column_2[16:23];
assign C24 = Column_2[24:31];

assign C31 = Column_3[0:7];
assign C32 = Column_3[8:15];
assign C33 = Column_3[16:23];
assign C34 = Column_3[24:31];

assign C41 = Column_4[0:7];
assign C42 = Column_4[8:15];
assign C43 = Column_4[16:23];
assign C44 = Column_4[24:31];

//

Multiply_By_14 A(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C11), .Read_Data(Q10));
Multiply_By_11 B(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C12), .Read_Data(Q11));
Multiply_By_13 C(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C13), .Read_Data(Q12));
Multiply_By_9 D(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C14), .Read_Data(Q13));

Multiply_By_14 E(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C12), .Read_Data(Q14));
Multiply_By_11 F(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C13), .Read_Data(Q15));
Multiply_By_13 G(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C14), .Read_Data(Q16));
Multiply_By_9 H(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C11), .Read_Data(Q17));

Multiply_By_14 I(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C13), .Read_Data(Q18));
Multiply_By_11 J(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C14), .Read_Data(Q19));
Multiply_By_13 K(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C11), .Read_Data(Q110));
Multiply_By_9 L(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C12), .Read_Data(Q111));

Multiply_By_14 M(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C14), .Read_Data(Q112));
Multiply_By_11 N(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C11), .Read_Data(Q113));
Multiply_By_13 O(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C12), .Read_Data(Q114));
Multiply_By_9 P(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C13), .Read_Data(Q115));

//

Multiply_By_14 Q(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C21), .Read_Data(Q20));
Multiply_By_11 R(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C22), .Read_Data(Q21));
Multiply_By_13 S(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C23), .Read_Data(Q22));
Multiply_By_9 T(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C24), .Read_Data(Q23));

Multiply_By_14 U(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C22), .Read_Data(Q24));
Multiply_By_11 V(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C23), .Read_Data(Q25));
Multiply_By_13 W(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C24), .Read_Data(Q26));
Multiply_By_9 X(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C21), .Read_Data(Q27));

Multiply_By_14 Y(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C23), .Read_Data(Q28));
Multiply_By_11 Z(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C24), .Read_Data(Q29));
Multiply_By_13 AA(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C21), .Read_Data(Q210));
Multiply_By_9 AB(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C22), .Read_Data(Q211));

Multiply_By_14 AC(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C24), .Read_Data(Q212));
Multiply_By_11 AD(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C21), .Read_Data(Q213));
Multiply_By_13 AE(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C22), .Read_Data(Q214));
Multiply_By_9 AF(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C23), .Read_Data(Q215));

//

Multiply_By_14 AG(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C31), .Read_Data(Q30));
Multiply_By_11 AH(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C32), .Read_Data(Q31));
Multiply_By_13 AI(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C33), .Read_Data(Q32));
Multiply_By_9 A1J(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C34), .Read_Data(Q33));

Multiply_By_14 AK(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C32), .Read_Data(Q34));
Multiply_By_11 AL(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C33), .Read_Data(Q35));
Multiply_By_13 AM(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C34), .Read_Data(Q36));
Multiply_By_9 AN(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C31), .Read_Data(Q37));

Multiply_By_14 AO(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C33), .Read_Data(Q38));
Multiply_By_11 AP(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C34), .Read_Data(Q39));
Multiply_By_13 AQ(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C31), .Read_Data(Q310));
Multiply_By_9 AR(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C32), .Read_Data(Q311));

Multiply_By_14 AS(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C34), .Read_Data(Q312));
Multiply_By_11 AT(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C31), .Read_Data(Q313));
Multiply_By_13 AU(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C32), .Read_Data(Q314));
Multiply_By_9 AV(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C33), .Read_Data(Q315));

//

Multiply_By_14 AW(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C41), .Read_Data(Q40));
Multiply_By_11 AX(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C42), .Read_Data(Q41));
Multiply_By_13 AY(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C43), .Read_Data(Q42));
Multiply_By_9 AZ(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C44), .Read_Data(Q43));

Multiply_By_14 BA(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C42), .Read_Data(Q44));
Multiply_By_11 BB(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C43), .Read_Data(Q45));
Multiply_By_13 BC(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C44), .Read_Data(Q46));
Multiply_By_9 BD(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C41), .Read_Data(Q47));

Multiply_By_14 BE(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C43), .Read_Data(Q48));
Multiply_By_11 BF(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C44), .Read_Data(Q49));
Multiply_By_13 BG(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C41), .Read_Data(Q410));
Multiply_By_9 BH(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C42), .Read_Data(Q411));

Multiply_By_14 BI(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C44), .Read_Data(Q412));
Multiply_By_11 BJ(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C41), .Read_Data(Q413));
Multiply_By_13 BK(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C42), .Read_Data(Q414));
Multiply_By_9 BL(.CLK(CLK), .Read_Enable(1'b1), .Read_Address(C43), .Read_Data(Q415));

//

assign OUTPUT[0:7] = (Q10 ^ Q11 ^ Q12 ^ Q13);
assign OUTPUT[8:15] = (Q14 ^ Q15 ^ Q16 ^ Q17);
assign OUTPUT[16:23] = (Q18 ^ Q19 ^ Q110 ^ Q111);
assign OUTPUT[24:31] = (Q112 ^ Q113 ^ Q114 ^ Q115);

assign OUTPUT[32:39] = (Q20 ^ Q21 ^ Q22 ^ Q23);
assign OUTPUT[40:47] = (Q24 ^ Q25 ^ Q26 ^ Q27);
assign OUTPUT[48:55] = (Q28 ^ Q29 ^ Q210 ^ Q211);
assign OUTPUT[56:63] = (Q212 ^ Q213 ^ Q214 ^ Q215);

assign OUTPUT[64:71] = (Q30 ^ Q31 ^ Q32 ^ Q33);
assign OUTPUT[72:79] = (Q34 ^ Q35 ^ Q36 ^ Q37);
assign OUTPUT[80:87] = (Q38 ^ Q39 ^ Q310 ^ Q311);
assign OUTPUT[88:95] = (Q312 ^ Q313 ^ Q314 ^ Q315);

assign OUTPUT[96:103] = (Q40 ^ Q41 ^ Q42 ^ Q43);
assign OUTPUT[104:111] = (Q44 ^ Q45 ^ Q46 ^ Q47);
assign OUTPUT[112:119] = (Q48 ^ Q49 ^ Q410 ^ Q411);
assign OUTPUT[120:127] = (Q412 ^ Q413 ^ Q414 ^ Q415);

endmodule

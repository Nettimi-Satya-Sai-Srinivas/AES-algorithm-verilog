module Input_Stage(
    input [0:127] INPUT,
    input [0:127] CIPHER_KEY,
    output [0:127] OUTPUT
    );

assign OUTPUT[0:7] = INPUT[0:7] ^ CIPHER_KEY[0:7];
assign OUTPUT[8:15] = INPUT[8:15] ^ CIPHER_KEY[8:15];
assign OUTPUT[16:23] = INPUT[16:23] ^ CIPHER_KEY[16:23];
assign OUTPUT[24:31] = INPUT[24:31] ^ CIPHER_KEY[24:31];

assign OUTPUT[32:39] = INPUT[32:39] ^ CIPHER_KEY[32:39];
assign OUTPUT[40:47] = INPUT[40:47] ^ CIPHER_KEY[40:47];
assign OUTPUT[48:55] = INPUT[48:55] ^ CIPHER_KEY[48:55];
assign OUTPUT[56:63] = INPUT[56:63] ^ CIPHER_KEY[56:63];

assign OUTPUT[64:71] = INPUT[64:71] ^ CIPHER_KEY[64:71];
assign OUTPUT[72:79] = INPUT[72:79] ^ CIPHER_KEY[72:79];
assign OUTPUT[80:87] = INPUT[80:87] ^ CIPHER_KEY[80:87];
assign OUTPUT[88:95] = INPUT[88:95] ^ CIPHER_KEY[88:95];

assign OUTPUT[96:103] = INPUT[96:103] ^ CIPHER_KEY[96:103];
assign OUTPUT[104:111] = INPUT[104:111] ^ CIPHER_KEY[104:111];
assign OUTPUT[112:119] = INPUT[112:119] ^ CIPHER_KEY[112:119];
assign OUTPUT[120:127] = INPUT[120:127] ^ CIPHER_KEY[120:127];

endmodule